-- synthesis library utils
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package fonts is
    type single_digit is array (0 to 7) of std_logic_vector(0 to 3);
    type digit_code is array(0 to 9) of single_digit;
    constant digits : digit_code := (
        ( -- 0
            "0000",
            "1110",
            "1010",
            "1010",
            "1010",
            "1110",
            "0000",
            "0000"
        ), -- 0
        ( -- 1
            "0000",
            "1000",
            "1000",
            "1000",
            "1000",
            "1000",
            "0000",
            "0000"
        ), -- 1
        ( -- 2
            "0000",
            "1110",
            "1000",
            "1110",
            "0010",
            "1110",
            "0000",
            "0000"
        ), -- 2
        ( -- 3
            "0000",
            "1110",
            "1000",
            "1100",
            "1000",
            "1110",
            "0000",
            "0000"
        ), -- 3
        ( -- 4
            "0000",
            "1010",
            "1010",
            "1110",
            "1000",
            "1000",
            "0000",
            "0000"
        ), -- 4
        ( -- 5
            "0000",
            "1110",
            "0010",
            "1110",
            "1000",
            "1110",
            "0000",
            "0000"
        ), -- 5
        ( -- 6
            "0000",
            "1110",
            "0010",
            "1110",
            "1010",
            "1110",
            "0000",
            "0000"
        ), -- 6
        ( -- 7
            "0000",
            "1110",
            "1000",
            "0100",
            "0010",
            "0010",
            "0000",
            "0000"
        ), -- 7
        ( -- 8
            "0000",
            "1110",
            "1010",
            "1110",
            "1010",
            "1110",
            "0000",
            "0000"
        ), -- 8
        ( -- 9
            "0000",
            "1110",
            "1010",
            "1110",
            "1000",
            "1110",
            "0000",
            "0000"
        ) -- 9
    );
end package fonts;
